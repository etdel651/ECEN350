module Decode24(out, in);
input [1:0] in;
output [3:0] out;

